//
`ifndef SV_STRING_PKG__SV
`define SV_STRING_PKG__SV

package sv_string_pkg;

    `include "sv_string_macros.svh"

    `include "sv_string_base.svh"

    `include "sv_string_function.svh"

endpackage

`endif
